--Instruction Memory and Instruction Decode
--
library ieee;
use ieee.std_logic_1164.all;

entity ARC_2 is
	port (PC_A: in std_logic_vector(31 downto 0);
			RS_A: out std_logic_vector(4 downto 0);		--5-bit RS output
			RT_A: out std_logic_vector(4 downto 0);		--5-bit RT output
			RD_A: out std_logic_vector(4 downto 0);		--5-bit RD output(R-Type only)
			IMM_A: out std_logic_vector(15 downto 0);	--5-bit IMM output(I-Type only)
			SHMT_A: out std_logic_vector(10 downto 6);	--5-bit Shift Amount (R-Type only)
			FUNCT_A: out std_logic_vector(5 downto 0);	--6-bit Function Code (R-Type only)
			TYPE_A: out std_logic_vector(1 downto 0));	--2-bit output to determine type: 00:R-Type, 01:J-Type, 10:I-Type, 11: error
end entity ARC_2;
	
architecture behave of ARC_2 is

signal TEMP_INST: std_logic_vector(31 downto 0);

component Instruction_Memory
	port (PC: in std_logic_vector(31 downto 0); 	--32-bit instruction
			INSTRUCTION: out std_logic_vector(31 downto 0)); --32-bit instruction(hardcoded in)
end component;

component Instruction_Decode 
	port (INST: in std_logic_vector(31 downto 0);    --32-bit instruction
			RS: out std_logic_vector(4 downto 0);		--5-bit RS output
			RT: out std_logic_vector(4 downto 0);		--5-bit RT output
			RD: out std_logic_vector(4 downto 0);		--5-bit RD output(R-Type only)
			IMM: out std_logic_vector(15 downto 0);		--5-bit IMM output(I-Type only)
			SHMT: out std_logic_vector(10 downto 6);	--5-bit Shift Amount (R-Type only)
			FUNCT: out std_logic_vector(5 downto 0);	--6-bit Function Code (R-Type only)
			TYPE_X: out std_logic_vector(1 downto 0));
			--TYPE: out std_logic_vector(1 downto 0);	--2-bit output to determine type: 00:R-Type, 01:J-Type, 10:I-Type, 11: error
end component;

begin

label1: Instruction_Memory port map(PC => PC_A, INSTRUCTION => TEMP_INST);
label2: Instruction_Decode port map(INST => TEMP_INST, RS => RS_A, RT => RT_A, RD => RD_A, IMM => IMM_A, SHMT => SHMT_A, FUNCT => FUNCT_A, TYPE_X => TYPE_A);
end architecture behave;	

